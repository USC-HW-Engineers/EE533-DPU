`timescale 1ns / 1ps
module gpu_top (
    input         clk,
    input         rst,
    input         run,
    input  [9:0]  thread_id,
    output        halted,
    output [9:0]  debug_pc,
    output [31:0] debug_ir,
    output [3:0]  debug_state
);

    // === Control Unit Signals ===
    wire [9:0]  pc;
    wire [4:0]  rf_rd_a, rf_rd_b, rf_rd_c, rf_wr_addr;
    wire        rf_we;
    wire [3:0]  alu_func;
    wire        tensor_start;
    wire [2:0]  tensor_op_mode;
    wire        tensor_relu_en;
    wire        dmem_we;
    wire [2:0]  wb_sel;
    wire [63:0] imm_out;
    wire [9:0]  dmem_addr;
    wire [3:0]  state;

    // === Instruction Memory ===
    wire [31:0] instruction;
    imem imem_inst (.clk(clk), .addr(pc), .data(instruction));

    // === Register File ===
    wire [63:0] rf_a, rf_b, rf_c;
    wire [63:0] rf_w_data;

    Register_file rf_inst (
        .clk(clk), .rst(rst), .we(rf_we),
        .w_addr(rf_wr_addr), .w_data(rf_w_data),
        .r_addr_a(rf_rd_a), .r_data_a(rf_a),
        .r_addr_b(rf_rd_b), .r_data_b(rf_b),
        .r_addr_c(rf_rd_c), .r_data_c(rf_c)
    );

    // === ALU ===
    wire [63:0] alu_result;
    alu alu_inst (
        .operand_a(rf_a), .operand_b(rf_b),
        .func(alu_func), .result(alu_result)
    );

    // === Tensor Unit ===
    wire [63:0] tensor_result;
    wire        tensor_done;
    tensor_unit tensor_inst (
        .clk(clk), .rst(rst), .start(tensor_start),
        .operand_a(rf_a), .operand_b(rf_b), .operand_c(rf_c),
        .op_mode(tensor_op_mode), .relu_en(tensor_relu_en),
        .result(tensor_result), .done(tensor_done)
    );

    // === Data Memory ===
    wire [63:0] dmem_rdata;
    dmem dmem_inst (
        .clk(clk), .we(dmem_we), .addr(dmem_addr),
        .w_data(rf_b), .r_data(dmem_rdata)
    );

    // === ReLU INT (per-lane max(0, x) on rf_a) ===
    wire [63:0] relu_int_result;
    assign relu_int_result[15:0]  = rf_a[15]  ? 16'b0 : rf_a[15:0];
    assign relu_int_result[31:16] = rf_a[31]  ? 16'b0 : rf_a[31:16];
    assign relu_int_result[47:32] = rf_a[47]  ? 16'b0 : rf_a[47:32];
    assign relu_int_result[63:48] = rf_a[63]  ? 16'b0 : rf_a[63:48];

    // === Writeback Mux ===
    reg [63:0] wb_data;
    always @(*) begin
        case (wb_sel)
            3'd0: wb_data = alu_result;
            3'd1: wb_data = tensor_result;
            3'd2: wb_data = dmem_rdata;
            3'd3: wb_data = imm_out;
            3'd4: wb_data = {54'b0, pc + 10'd1};
            3'd5: wb_data = imm_out;
            3'd6: wb_data = relu_int_result;
            default: wb_data = 64'b0;
        endcase
    end

    assign rf_w_data = wb_data;

    // === Control Unit ===
    control_unit ctrl_inst (
        .clk(clk), .rst(rst), .run(run),
        .instruction(instruction), .tensor_done(tensor_done),
        .thread_id(thread_id),
        .cmp_a(rf_a), .cmp_b(rf_b),
        .pc(pc),
        .rf_rd_a(rf_rd_a), .rf_rd_b(rf_rd_b), .rf_rd_c(rf_rd_c),
        .rf_wr_addr(rf_wr_addr), .rf_we(rf_we),
        .alu_func(alu_func),
        .tensor_start(tensor_start), .tensor_op_mode(tensor_op_mode),
        .tensor_relu_en(tensor_relu_en),
        .dmem_we(dmem_we), .wb_sel(wb_sel),
        .imm_out(imm_out), .dmem_addr(dmem_addr),
        .halted(halted), .state(state)
    );

    // === Debug Outputs ===
    assign debug_pc    = pc;
    assign debug_ir    = instruction;
    assign debug_state = state;

endmodule
